`define         ADR_WIDTH           32
`define         PCADR_WIDTH     16
`define         DATA_WIDTH      32
`define         RST_VALID       1'b1
`define         VALID_EN        1'b1
`define         ADDR_WIDTH      32
`define         DATA_WIDTH      32
`define         REG_WRITE       1'b1
`define         ALUADD          4'b0010
`define         ALUADDU         4'b0000
`define         ALUSUB          4'b0011
`define         ALUAND          4'b0100
`define         ALUOR           4'b0101
`define         ALUXOR          4'b0110
`define         ALUNOR          4'b0111
`define         ALUSLT          4'b1011
`define         ALUSLTU         4'b1010
`define         ALUEQU          4'b0001
`define         ALUNEQ          4'b1100
`define         ALUSLL          4'b1000
`define         ALUSRA          4'b1001
`define         ALUSRL          4'b1101